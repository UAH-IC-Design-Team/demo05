`default_nettype none
`timescale 10ns/1ns

module clk_div(
);

endmodule
